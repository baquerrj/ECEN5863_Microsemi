library IEEE;
use IEEE.std_logic_1164.all;

entity MSS_APB is

  generic
  (
    ACT_CONFIG : integer := 0;
    ACT_FCLK   : integer := 0;
    ACT_DIE    : string := "";
    ACT_PKG    : string := ""
  );

  port
  (
    ABPS0            : in  std_logic;
    ABPS1            : in  std_logic;
    ABPS10           : in  std_logic;
    ABPS11           : in  std_logic;
    ABPS2            : in  std_logic;
    ABPS3            : in  std_logic;
    ABPS4            : in  std_logic;
    ABPS5            : in  std_logic;
    ABPS6            : in  std_logic;
    ABPS7            : in  std_logic;
    ABPS8            : in  std_logic;
    ABPS9            : in  std_logic;
    ACEFLAGS         : out std_logic_vector(31 downto 0);
    ADC0             : in  std_logic;
    ADC1             : in  std_logic;
    ADC10            : in  std_logic;
    ADC11            : in  std_logic;
    ADC2             : in  std_logic;
    ADC3             : in  std_logic;
    ADC4             : in  std_logic;
    ADC5             : in  std_logic;
    ADC6             : in  std_logic;
    ADC7             : in  std_logic;
    ADC8             : in  std_logic;
    ADC9             : in  std_logic;
    CALIBIN          : in  std_logic;
    CALIBOUT         : out std_logic;
    CM0              : in  std_logic;
    CM1              : in  std_logic;
    CM2              : in  std_logic;
    CM3              : in  std_logic;
    CM4              : in  std_logic;
    CM5              : in  std_logic;
    CMP0             : out std_logic;
    CMP1             : out std_logic;
    CMP10            : out std_logic;
    CMP11            : out std_logic;
    CMP2             : out std_logic;
    CMP3             : out std_logic;
    CMP4             : out std_logic;
    CMP5             : out std_logic;
    CMP6             : out std_logic;
    CMP7             : out std_logic;
    CMP8             : out std_logic;
    CMP9             : out std_logic;
    DEEPSLEEP        : out std_logic;
    DMAREADY         : in  std_logic_vector(1 downto 0);
    EMCAB            : out std_logic_vector(25 downto 0);
    EMCBYTEN         : out std_logic_vector(1 downto 0);
    EMCCLK           : out std_logic;
    EMCCLKRTN        : in  std_logic;
    EMCCS0n          : out std_logic;
    EMCCS1n          : out std_logic;
    EMCDBOE          : out std_logic;
    EMCOEN0n         : out std_logic;
    EMCOEN1n         : out std_logic;
    EMCRDB           : in  std_logic_vector(15 downto 0);
    EMCRWn           : out std_logic;
    EMCWDB           : out std_logic_vector(15 downto 0);
    F2MRESETn        : in  std_logic;
    FABACETRIG       : in  std_logic;
    FABINT           : in  std_logic;
    FABPADDR         : in  std_logic_vector(31 downto 0);
    FABPENABLE       : in  std_logic;
    FABPRDATA        : out std_logic_vector(31 downto 0);
    FABPREADY        : out std_logic;
    FABPSEL          : in  std_logic;
    FABPSLVERR       : out std_logic;
    FABPWDATA        : in  std_logic_vector(31 downto 0);
    FABPWRITE        : in  std_logic;
    FABSDD0CLK       : in  std_logic;
    FABSDD0D         : in  std_logic;
    FABSDD1CLK       : in  std_logic;
    FABSDD1D         : in  std_logic;
    FABSDD2CLK       : in  std_logic;
    FABSDD2D         : in  std_logic;
    FCLK             : in  std_logic;
    GNDTM0           : in  std_logic;
    GNDTM1           : in  std_logic;
    GNDTM2           : in  std_logic;
    GNDVAREF         : in  std_logic;
    GPI              : in  std_logic_vector(31 downto 0);
    GPO              : out std_logic_vector(31 downto 0);
    GPOE             : out std_logic_vector(31 downto 0);
    I2C0BCLK         : in  std_logic;
    I2C0SCLI         : in  std_logic;
    I2C0SCLO         : out std_logic;
    I2C0SDAI         : in  std_logic;
    I2C0SDAO         : out std_logic;
    I2C0SMBALERTNI   : in  std_logic;
    I2C0SMBALERTNO   : out std_logic;
    I2C0SMBUSNI      : in  std_logic;
    I2C0SMBUSNO      : out std_logic;
    I2C1BCLK         : in  std_logic;
    I2C1SCLI         : in  std_logic;
    I2C1SCLO         : out std_logic;
    I2C1SDAI         : in  std_logic;
    I2C1SDAO         : out std_logic;
    I2C1SMBALERTNI   : in  std_logic;
    I2C1SMBALERTNO   : out std_logic;
    I2C1SMBUSNI      : in  std_logic;
    I2C1SMBUSNO      : out std_logic;
    LVTTL0           : out std_logic;
    LVTTL0EN         : in  std_logic;
    LVTTL1           : out std_logic;
    LVTTL10          : out std_logic;
    LVTTL10EN        : in  std_logic;
    LVTTL11          : out std_logic;
    LVTTL11EN        : in  std_logic;
    LVTTL1EN         : in  std_logic;
    LVTTL2           : out std_logic;
    LVTTL2EN         : in  std_logic;
    LVTTL3           : out std_logic;
    LVTTL3EN         : in  std_logic;
    LVTTL4           : out std_logic;
    LVTTL4EN         : in  std_logic;
    LVTTL5           : out std_logic;
    LVTTL5EN         : in  std_logic;
    LVTTL6           : out std_logic;
    LVTTL6EN         : in  std_logic;
    LVTTL7           : out std_logic;
    LVTTL7EN         : in  std_logic;
    LVTTL8           : out std_logic;
    LVTTL8EN         : in  std_logic;
    LVTTL9           : out std_logic;
    LVTTL9EN         : in  std_logic;
    M2FRESETn        : out std_logic;
    MACCLK           : in  std_logic;
    MACCLKCCC        : in  std_logic;
    MACCRSDV         : in  std_logic;
    MACF2MCRSDV      : in  std_logic;
    MACF2MMDI        : in  std_logic;
    MACF2MRXD        : in  std_logic_vector(1 downto 0);
    MACF2MRXER       : in  std_logic;
    MACM2FMDC        : out std_logic;
    MACM2FMDEN       : out std_logic;
    MACM2FMDO        : out std_logic;
    MACM2FTXD        : out std_logic_vector(1 downto 0);
    MACM2FTXEN       : out std_logic;
    MACMDC           : out std_logic;
    MACMDEN          : out std_logic;
    MACMDI           : in  std_logic;
    MACMDO           : out std_logic;
    MACRXD           : in  std_logic_vector(1 downto 0);
    MACRXER          : in  std_logic;
    MACTXD           : out std_logic_vector(1 downto 0);
    MACTXEN          : out std_logic;
    MSSINT           : out std_logic_vector(7 downto 0);
    MSSPADDR         : out std_logic_vector(19 downto 0);
    MSSPENABLE       : out std_logic;
    MSSPRDATA        : in  std_logic_vector(31 downto 0);
    MSSPREADY        : in  std_logic;
    MSSPSEL          : out std_logic;
    MSSPSLVERR       : in  std_logic;
    MSSPWDATA        : out std_logic_vector(31 downto 0);
    MSSPWRITE        : out std_logic;
    MSSRESETn        : in  std_logic;
    PLLLOCK          : in  std_logic;
    PUFABn           : out std_logic;
    PUn              : in  std_logic;
    RCOSC            : in  std_logic;
    RXEV             : in  std_logic;
    SDD0             : out std_logic;
    SDD1             : out std_logic;
    SDD2             : out std_logic;
    SLEEP            : out std_logic;
    SPI0CLKI         : in  std_logic;
    SPI0CLKO         : out std_logic;
    SPI0DI           : in  std_logic;
    SPI0DO           : out std_logic;
    SPI0DOE          : out std_logic;
    SPI0MODE         : out std_logic;
    SPI0SSI          : in  std_logic;
    SPI0SSO          : out std_logic_vector(7 downto 0);
    SPI1CLKI         : in  std_logic;
    SPI1CLKO         : out std_logic;
    SPI1DI           : in  std_logic;
    SPI1DO           : out std_logic;
    SPI1DOE          : out std_logic;
    SPI1MODE         : out std_logic;
    SPI1SSI          : in  std_logic;
    SPI1SSO          : out std_logic_vector(7 downto 0);
    SYNCCLKFDBK      : in  std_logic;
    TM0              : in  std_logic;
    TM1              : in  std_logic;
    TM2              : in  std_logic;
    TM3              : in  std_logic;
    TM4              : in  std_logic;
    TM5              : in  std_logic;
    TXEV             : out std_logic;
    UART0CTSn        : in  std_logic;
    UART0DCDn        : in  std_logic;
    UART0DSRn        : in  std_logic;
    UART0DTRn        : out std_logic;
    UART0RIn         : in  std_logic;
    UART0RTSn        : out std_logic;
    UART0RXD         : in  std_logic;
    UART0TXD         : out std_logic;
    UART1CTSn        : in  std_logic;
    UART1DCDn        : in  std_logic;
    UART1DSRn        : in  std_logic;
    UART1DTRn        : out std_logic;
    UART1RIn         : in  std_logic;
    UART1RTSn        : out std_logic;
    UART1RXD         : in  std_logic;
    UART1TXD         : out std_logic;
    VAREF0           : in  std_logic;
    VAREF1           : in  std_logic;
    VAREF2           : in  std_logic;
    VAREFOUT         : out std_logic;
    VCC15GOOD        : out std_logic;
    VCC33GOOD        : out std_logic;
    VRON             : in  std_logic;
    WDINT            : out std_logic
  );

end MSS_APB;

architecture DEF_ARCH of MSS_APB is

    attribute syn_black_box : boolean;
    attribute syn_black_box of DEF_ARCH : architecture is true;
    attribute syn_tco1 : string;
    attribute syn_tco1 of DEF_ARCH : architecture is "FCLK->ACEFLAGS[31:0]=5.641";
    attribute syn_tco2 : string;
    attribute syn_tco2 of DEF_ARCH : architecture is "FCLK->DEEPSLEEP=3.492";
    attribute syn_tsu1 : string;
    attribute syn_tsu1 of DEF_ARCH : architecture is "DMAREADY[1:0]->FCLK=1.468";
    attribute syn_tco3 : string;
    attribute syn_tco3 of DEF_ARCH : architecture is "FCLK->EMCAB[25:0]=2.672";
    attribute syn_tco4 : string;
    attribute syn_tco4 of DEF_ARCH : architecture is "FCLK->EMCBYTEN[1:0]=4.324";
    attribute syn_tco5 : string;
    attribute syn_tco5 of DEF_ARCH : architecture is "FCLK->EMCCS0n=4.522";
    attribute syn_tco6 : string;
    attribute syn_tco6 of DEF_ARCH : architecture is "FCLK->EMCCS1n=4.554";
    attribute syn_tco7 : string;
    attribute syn_tco7 of DEF_ARCH : architecture is "FCLK->EMCDBOE=2.672";
    attribute syn_tco8 : string;
    attribute syn_tco8 of DEF_ARCH : architecture is "FCLK->EMCOEN0n=4.303";
    attribute syn_tco9 : string;
    attribute syn_tco9 of DEF_ARCH : architecture is "FCLK->EMCOEN1n=4.314";
    attribute syn_tsu2 : string;
    attribute syn_tsu2 of DEF_ARCH : architecture is "EMCRDB[15:0]->EMCCLKRTN=0.003";
    attribute syn_tco10 : string;
    attribute syn_tco10 of DEF_ARCH : architecture is "FCLK->EMCRWn=2.924";
    attribute syn_tco11 : string;
    attribute syn_tco11 of DEF_ARCH : architecture is "FCLK->EMCWDB[15:0]=6.91";
    attribute syn_tsu3 : string;
    attribute syn_tsu3 of DEF_ARCH : architecture is "FABACETRIG->FCLK=0";
    attribute syn_tsu4 : string;
    attribute syn_tsu4 of DEF_ARCH : architecture is "FABINT->FCLK=0.321";
    attribute syn_tsu5 : string;
    attribute syn_tsu5 of DEF_ARCH : architecture is "FABPADDR[31:0]->FCLK=0";
    attribute syn_tsu6 : string;
    attribute syn_tsu6 of DEF_ARCH : architecture is "FABPENABLE->FCLK=0";
    attribute syn_tco12 : string;
    attribute syn_tco12 of DEF_ARCH : architecture is "FCLK->FABPRDATA[31:0]=3.926";
    attribute syn_tco13 : string;
    attribute syn_tco13 of DEF_ARCH : architecture is "FCLK->FABPREADY=2.712";
    attribute syn_tsu7 : string;
    attribute syn_tsu7 of DEF_ARCH : architecture is "FABPSEL->FCLK=0";
    attribute syn_tco14 : string;
    attribute syn_tco14 of DEF_ARCH : architecture is "FCLK->FABPSLVERR=2.859";
    attribute syn_tsu8 : string;
    attribute syn_tsu8 of DEF_ARCH : architecture is "FABPWDATA[31:0]->FCLK=0";
    attribute syn_tsu9 : string;
    attribute syn_tsu9 of DEF_ARCH : architecture is "FABPWRITE->FCLK=0";
    attribute syn_tsu10 : string;
    attribute syn_tsu10 of DEF_ARCH : architecture is "GPI[31:0]->FCLK=0.516";
    attribute syn_tco15 : string;
    attribute syn_tco15 of DEF_ARCH : architecture is "FCLK->GPO[31:0]=4.132";
    attribute syn_tco16 : string;
    attribute syn_tco16 of DEF_ARCH : architecture is "FCLK->GPOE[31:0]=3.908";
    attribute syn_tsu11 : string;
    attribute syn_tsu11 of DEF_ARCH : architecture is "I2C0BCLK->FCLK=0";
    attribute syn_tsu12 : string;
    attribute syn_tsu12 of DEF_ARCH : architecture is "I2C0SCLI->FCLK=0";
    attribute syn_tco17 : string;
    attribute syn_tco17 of DEF_ARCH : architecture is "FCLK->I2C0SCLO=3.465";
    attribute syn_tsu13 : string;
    attribute syn_tsu13 of DEF_ARCH : architecture is "I2C0SDAI->FCLK=0";
    attribute syn_tco18 : string;
    attribute syn_tco18 of DEF_ARCH : architecture is "FCLK->I2C0SDAO=3.368";
    attribute syn_tsu14 : string;
    attribute syn_tsu14 of DEF_ARCH : architecture is "I2C0SMBALERTNI->FCLK=0";
    attribute syn_tco19 : string;
    attribute syn_tco19 of DEF_ARCH : architecture is "FCLK->I2C0SMBALERTNO=2.855";
    attribute syn_tsu15 : string;
    attribute syn_tsu15 of DEF_ARCH : architecture is "I2C0SMBUSNI->FCLK=0";
    attribute syn_tco20 : string;
    attribute syn_tco20 of DEF_ARCH : architecture is "FCLK->I2C0SMBUSNO=2.916";
    attribute syn_tsu16 : string;
    attribute syn_tsu16 of DEF_ARCH : architecture is "I2C1BCLK->FCLK=0";
    attribute syn_tsu17 : string;
    attribute syn_tsu17 of DEF_ARCH : architecture is "I2C1SCLI->FCLK=0";
    attribute syn_tco21 : string;
    attribute syn_tco21 of DEF_ARCH : architecture is "FCLK->I2C1SCLO=3.762";
    attribute syn_tsu18 : string;
    attribute syn_tsu18 of DEF_ARCH : architecture is "I2C1SDAI->FCLK=0.045";
    attribute syn_tco22 : string;
    attribute syn_tco22 of DEF_ARCH : architecture is "FCLK->I2C1SDAO=3.712";
    attribute syn_tsu19 : string;
    attribute syn_tsu19 of DEF_ARCH : architecture is "I2C1SMBALERTNI->FCLK=0";
    attribute syn_tco23 : string;
    attribute syn_tco23 of DEF_ARCH : architecture is "FCLK->I2C1SMBALERTNO=2.5";
    attribute syn_tsu20 : string;
    attribute syn_tsu20 of DEF_ARCH : architecture is "I2C1SMBUSNI->FCLK=0";
    attribute syn_tco24 : string;
    attribute syn_tco24 of DEF_ARCH : architecture is "FCLK->I2C1SMBUSNO=2.501";
    attribute syn_tco25 : string;
    attribute syn_tco25 of DEF_ARCH : architecture is "FCLK->M2FRESETn=2.957";
    attribute syn_tsu21 : string;
    attribute syn_tsu21 of DEF_ARCH : architecture is "MACCRSDV->MACCLK=0";
    attribute syn_tsu22 : string;
    attribute syn_tsu22 of DEF_ARCH : architecture is "MACCRSDV->MACCLKCCC=0";
    attribute syn_tsu23 : string;
    attribute syn_tsu23 of DEF_ARCH : architecture is "MACF2MCRSDV->MACCLK=0";
    attribute syn_tsu24 : string;
    attribute syn_tsu24 of DEF_ARCH : architecture is "MACF2MCRSDV->MACCLKCCC=0";
    attribute syn_tsu25 : string;
    attribute syn_tsu25 of DEF_ARCH : architecture is "MACF2MMDI->FCLK=0";
    attribute syn_tsu26 : string;
    attribute syn_tsu26 of DEF_ARCH : architecture is "MACF2MRXD[1:0]->MACCLK=0";
    attribute syn_tsu27 : string;
    attribute syn_tsu27 of DEF_ARCH : architecture is "MACF2MRXD[1:0]->MACCLKCCC=0";
    attribute syn_tsu28 : string;
    attribute syn_tsu28 of DEF_ARCH : architecture is "MACF2MRXER->MACCLK=0";
    attribute syn_tsu29 : string;
    attribute syn_tsu29 of DEF_ARCH : architecture is "MACF2MRXER->MACCLKCCC=0";
    attribute syn_tco26 : string;
    attribute syn_tco26 of DEF_ARCH : architecture is "FCLK->MACM2FMDC=3.861";
    attribute syn_tco27 : string;
    attribute syn_tco27 of DEF_ARCH : architecture is "FCLK->MACM2FMDEN=4.061";
    attribute syn_tco28 : string;
    attribute syn_tco28 of DEF_ARCH : architecture is "FCLK->MACM2FMDO=4.261";
    attribute syn_tco29 : string;
    attribute syn_tco29 of DEF_ARCH : architecture is "FCLK->MACM2FTXD[1:0]=3.912";
    attribute syn_tco30 : string;
    attribute syn_tco30 of DEF_ARCH : architecture is "MACCLK->MACM2FTXD[1:0]=2.855";
    attribute syn_tco31 : string;
    attribute syn_tco31 of DEF_ARCH : architecture is "FCLK->MACM2FTXEN=4.167";
    attribute syn_tco32 : string;
    attribute syn_tco32 of DEF_ARCH : architecture is "MACCLK->MACM2FTXEN=2.843";
    attribute syn_tco33 : string;
    attribute syn_tco33 of DEF_ARCH : architecture is "FCLK->MACMDC=3.198";
    attribute syn_tco34 : string;
    attribute syn_tco34 of DEF_ARCH : architecture is "FCLK->MACMDEN=3.664";
    attribute syn_tsu30 : string;
    attribute syn_tsu30 of DEF_ARCH : architecture is "MACMDI->FCLK=0";
    attribute syn_tco35 : string;
    attribute syn_tco35 of DEF_ARCH : architecture is "FCLK->MACMDO=3.524";
    attribute syn_tsu31 : string;
    attribute syn_tsu31 of DEF_ARCH : architecture is "MACRXD[1:0]->MACCLK=0";
    attribute syn_tsu32 : string;
    attribute syn_tsu32 of DEF_ARCH : architecture is "MACRXD[1:0]->MACCLKCCC=0";
    attribute syn_tsu33 : string;
    attribute syn_tsu33 of DEF_ARCH : architecture is "MACRXER->MACCLK=0";
    attribute syn_tsu34 : string;
    attribute syn_tsu34 of DEF_ARCH : architecture is "MACRXER->MACCLKCCC=0";
    attribute syn_tco36 : string;
    attribute syn_tco36 of DEF_ARCH : architecture is "FCLK->MACTXD[1:0]=3.24";
    attribute syn_tco37 : string;
    attribute syn_tco37 of DEF_ARCH : architecture is "MACCLK->MACTXD[1:0]=2.596";
    attribute syn_tco38 : string;
    attribute syn_tco38 of DEF_ARCH : architecture is "FCLK->MACTXEN=3.601";
    attribute syn_tco39 : string;
    attribute syn_tco39 of DEF_ARCH : architecture is "MACCLK->MACTXEN=2.745";
    attribute syn_tco40 : string;
    attribute syn_tco40 of DEF_ARCH : architecture is "FCLK->MSSINT[7:0]=5.637";
    attribute syn_tco41 : string;
    attribute syn_tco41 of DEF_ARCH : architecture is "FCLK->MSSPADDR[19:0]=2.679";
    attribute syn_tco42 : string;
    attribute syn_tco42 of DEF_ARCH : architecture is "FCLK->MSSPENABLE=2.474";
    attribute syn_tsu35 : string;
    attribute syn_tsu35 of DEF_ARCH : architecture is "MSSPRDATA[31:0]->FCLK=0";
    attribute syn_tsu36 : string;
    attribute syn_tsu36 of DEF_ARCH : architecture is "MSSPREADY->FCLK=0";
    attribute syn_tco43 : string;
    attribute syn_tco43 of DEF_ARCH : architecture is "FCLK->MSSPSEL=2.49";
    attribute syn_tsu37 : string;
    attribute syn_tsu37 of DEF_ARCH : architecture is "MSSPSLVERR->FCLK=0";
    attribute syn_tco44 : string;
    attribute syn_tco44 of DEF_ARCH : architecture is "FCLK->MSSPWDATA[31:0]=2.71";
    attribute syn_tco45 : string;
    attribute syn_tco45 of DEF_ARCH : architecture is "FCLK->MSSPWRITE=2.456";
    attribute syn_tsu38 : string;
    attribute syn_tsu38 of DEF_ARCH : architecture is "MSSRESETn->FCLK=0";
    attribute syn_tsu39 : string;
    attribute syn_tsu39 of DEF_ARCH : architecture is "PUn->FCLK=0";
    attribute syn_tsu40 : string;
    attribute syn_tsu40 of DEF_ARCH : architecture is "RXEV->FCLK=0";
    attribute syn_tco46 : string;
    attribute syn_tco46 of DEF_ARCH : architecture is "FCLK->SLEEP=3.304";
    attribute syn_tsu41 : string;
    attribute syn_tsu41 of DEF_ARCH : architecture is "SPI0CLKI->FCLK=0";
    attribute syn_tco47 : string;
    attribute syn_tco47 of DEF_ARCH : architecture is "FCLK->SPI0CLKO=3.407";
    attribute syn_tsu42 : string;
    attribute syn_tsu42 of DEF_ARCH : architecture is "SPI0DI->FCLK=0";
    attribute syn_tco48 : string;
    attribute syn_tco48 of DEF_ARCH : architecture is "FCLK->SPI0DO=4.35";
    attribute syn_tco49 : string;
    attribute syn_tco49 of DEF_ARCH : architecture is "FCLK->SPI0DOE=4.947";
    attribute syn_tco50 : string;
    attribute syn_tco50 of DEF_ARCH : architecture is "FCLK->SPI0MODE=3.423";
    attribute syn_tsu43 : string;
    attribute syn_tsu43 of DEF_ARCH : architecture is "SPI0SSI->FCLK=0.858";
    attribute syn_tco51 : string;
    attribute syn_tco51 of DEF_ARCH : architecture is "FCLK->SPI0SSO[7:0]=4.117";
    attribute syn_tsu44 : string;
    attribute syn_tsu44 of DEF_ARCH : architecture is "SPI1CLKI->FCLK=0";
    attribute syn_tco52 : string;
    attribute syn_tco52 of DEF_ARCH : architecture is "FCLK->SPI1CLKO=3.548";
    attribute syn_tsu45 : string;
    attribute syn_tsu45 of DEF_ARCH : architecture is "SPI1DI->FCLK=0";
    attribute syn_tco53 : string;
    attribute syn_tco53 of DEF_ARCH : architecture is "FCLK->SPI1DO=4.643";
    attribute syn_tco54 : string;
    attribute syn_tco54 of DEF_ARCH : architecture is "FCLK->SPI1DOE=4.318";
    attribute syn_tco55 : string;
    attribute syn_tco55 of DEF_ARCH : architecture is "FCLK->SPI1MODE=4.136";
    attribute syn_tsu46 : string;
    attribute syn_tsu46 of DEF_ARCH : architecture is "SPI1SSI->FCLK=0.271";
    attribute syn_tco56 : string;
    attribute syn_tco56 of DEF_ARCH : architecture is "FCLK->SPI1SSO[7:0]=4.904";
    attribute syn_tco57 : string;
    attribute syn_tco57 of DEF_ARCH : architecture is "FCLK->TXEV=4.597";
    attribute syn_tsu47 : string;
    attribute syn_tsu47 of DEF_ARCH : architecture is "UART0CTSn->FCLK=0";
    attribute syn_tsu48 : string;
    attribute syn_tsu48 of DEF_ARCH : architecture is "UART0DCDn->FCLK=0";
    attribute syn_tsu49 : string;
    attribute syn_tsu49 of DEF_ARCH : architecture is "UART0DSRn->FCLK=0";
    attribute syn_tco58 : string;
    attribute syn_tco58 of DEF_ARCH : architecture is "FCLK->UART0DTRn=3.299";
    attribute syn_tsu50 : string;
    attribute syn_tsu50 of DEF_ARCH : architecture is "UART0RIn->FCLK=0";
    attribute syn_tco59 : string;
    attribute syn_tco59 of DEF_ARCH : architecture is "FCLK->UART0RTSn=3.349";
    attribute syn_tsu51 : string;
    attribute syn_tsu51 of DEF_ARCH : architecture is "UART0RXD->FCLK=0.076";
    attribute syn_tco60 : string;
    attribute syn_tco60 of DEF_ARCH : architecture is "FCLK->UART0TXD=3.571";
    attribute syn_tsu52 : string;
    attribute syn_tsu52 of DEF_ARCH : architecture is "UART1CTSn->FCLK=0";
    attribute syn_tsu53 : string;
    attribute syn_tsu53 of DEF_ARCH : architecture is "UART1DCDn->FCLK=0";
    attribute syn_tsu54 : string;
    attribute syn_tsu54 of DEF_ARCH : architecture is "UART1DSRn->FCLK=0";
    attribute syn_tco61 : string;
    attribute syn_tco61 of DEF_ARCH : architecture is "FCLK->UART1DTRn=3.407";
    attribute syn_tsu55 : string;
    attribute syn_tsu55 of DEF_ARCH : architecture is "UART1RIn->FCLK=0";
    attribute syn_tco62 : string;
    attribute syn_tco62 of DEF_ARCH : architecture is "FCLK->UART1RTSn=3.714";
    attribute syn_tsu56 : string;
    attribute syn_tsu56 of DEF_ARCH : architecture is "UART1RXD->FCLK=0";
    attribute syn_tco63 : string;
    attribute syn_tco63 of DEF_ARCH : architecture is "FCLK->UART1TXD=3.585";
    attribute syn_tco64 : string;
    attribute syn_tco64 of DEF_ARCH : architecture is "FCLK->WDINT=2.749";

begin
end DEF_ARCH;
